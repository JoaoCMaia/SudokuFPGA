
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Cronometer is
     PORT (
         clk : in  STD_LOGIC;
         rst: in STD_LOGIC;         
         colorOutClock : out  STD_LOGIC_VECTOR(11 DOWNTO 0);
         current_x: in STD_LOGIC_VECTOR(9 downto 0);
         current_y: in STD_LOGIC_VECTOR(9 downto 0);
         second:out std_logic_vector(3 downto 0);
         finish: in std_logic
         
 );
end Cronometer;

architecture Behavioral of Cronometer is
 TYPE digit18x24 IS ARRAY (1 TO 24, 1 TO 18) OF STD_LOGIC;
  CONSTANT zero: digit18x24 :=(
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')); 
 CONSTANT one: digit18x24 := (
	    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0'),
        ('0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
    CONSTANT two: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));    
    CONSTANT three: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
    CONSTANT four: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),        
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')); 
    CONSTANT five: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
    CONSTANT six: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
    CONSTANT seven: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
    CONSTANT eight: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));  
    CONSTANT nine: digit18x24 := (
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
        ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')); 
         TYPE digit46x14 IS ARRAY (1 TO 14, 1 TO 46) OF STD_LOGIC;
         CONSTANT Win: digit46x14 :=(
        ('1','1','1','1','1','1','0','0','0','0','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1'),
        ('0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1'),
        ('0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0'),
        ('0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','1','1','0','0','0','0','0','1','0','0'),
        ('0','0','0','1','1','0','0','0','1','0','0','1','0','0','0','0','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','1','1','1','0','0','0','0','1','0','0'),
        ('0','0','0','1','1','0','0','0','1','0','0','1','1','0','0','0','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','1','1','0','0','0','0','1','0','0'),
        ('0','0','0','1','1','0','0','0','1','0','0','1','1','0','0','0','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','1','1','0','0','0','1','0','0'),
        ('0','0','0','1','1','1','0','1','0','0','0','1','1','0','0','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','1','1','1','0','0','1','0','0'),
        ('0','0','0','0','1','1','0','1','0','0','0','0','1','1','0','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','0','1','1','0','0','1','0','0'),
        ('0','0','0','0','1','1','0','1','0','0','0','0','1','1','0','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','1','1','0','1','0','0'),
        ('0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','1','0','0'),
        ('0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','1','0','0'),
        ('0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0'),
        ('0','0','0','0','0','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','0','0'));    
        CONSTANT MAX_WIDTH: natural :=27;
        constant DIGITHIGH: natural:=23;
        constant DIGITLENGHT: natural:=17;
        constant FINALHIGH: natural :=(231);
        constant all_ones : std_logic_vector (MAX_WIDTH-1 downto 0) := "101111101011110000100000000";
        signal counter : std_logic_vector (MAX_WIDTH-1 downto 0) := (others =>'0');
        signal ctick: std_logic :='0';
        signal unidade, dezenas, centenas, milhar : std_logic_vector(3 downto 0) :=(others=>'0');
        signal colorOut : STD_LOGIC_VECTOR(11 DOWNTO 0);
        
        ---Function construction:----------------
     FUNCTION bcd_to_digit6x8 (SIGNAL input: std_logic_vector(3 downto 0)) RETURN digit18x24 IS
     BEGIN
         CASE input is
             WHEN "0000" => return zero;
             WHEN "0001" => return one;
             WHEN "0010" => return two;
             WHEN "0011" => return three;
             WHEN "0100" => return four;
             WHEN "0101" => return five;
             WHEN "0110" => return six;
             WHEN "0111" => return seven;
             WHEN "1000" => return eight;
             WHEN "1001" => return nine;
             when others => return zero;
         END CASE;
     END bcd_to_digit6x8;
    -------------------------------------------
    
begin
    colorOutClock<=colorOut;
    
    process(clk,counter)
    begin
        if rising_edge (clk)then
            counter <= counter + 1;
            if counter = all_ones then
                ctick <= '1';
                counter <=(others=>'0');
            else
                ctick <= '0';
            end if;
        end if;    
    end process;
    second<=unidade;
    process(clk,ctick, unidade, dezenas,centenas,milhar, finish)
       begin
        if (rising_edge(clk) and finish='0')then
           if(rst='1')then
                unidade<=(others=>'0');
                dezenas<=(others=>'0');
                centenas<=(others=>'0');
                milhar<=(others=>'0');
           else 
               if(ctick='1')then    
                   unidade<= unidade + 1;
                        if unidade = "1001" then
                            dezenas<= dezenas +1;
                            unidade<=(others=>'0');
                            if dezenas = "1001" then
                               centenas<= centenas +1;
                               dezenas<=(others=>'0');
                                if centenas = "1001" then
                                   milhar<= milhar +1;
                                   centenas<=(others=>'0');
                                end if;
                             end if;
                        end if;
                end if;    
             end if;           
        end if;          
    end process;

    process(finish, unidade, dezenas,centenas,milhar,counter, current_x, current_y) 
    begin
        colorOut<= (others=>'0');
        if(finish='0')then
            IF(current_x >= x"236" AND current_x < (x"236"+ DIGITLENGHT) AND current_y >=  x"01" AND current_y < (x"01" + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(milhar)(to_Integer(UNSIGNED(current_y- x"01")),to_Integer(UNSIGNED(current_x- x"236"))));
            elsIF(current_x >= x"249" AND current_x < (x"249"+ DIGITLENGHT) AND current_y >=  x"01" AND current_y < (x"01" + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(centenas)(to_Integer(UNSIGNED(current_y- x"01")),to_Integer(UNSIGNED(current_x- x"249"))));
            elsIF(current_x >= x"25C" AND current_x < (x"25C"+ DIGITLENGHT) AND current_y >=  x"01" AND current_y < (x"01" + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(dezenas)(to_Integer(UNSIGNED(current_y- x"01")),to_Integer(UNSIGNED(current_x- x"25C"))));
            elsIF(current_x >= x"26F" AND current_x < (x"26F"+ DIGITLENGHT) AND current_y >=  x"01" AND current_y < (x"01" + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(unidade)(to_Integer(UNSIGNED(current_y- x"01")),to_Integer(UNSIGNED(current_x- x"26F"))));
            end if;
        else
            IF(current_x >= x"10E" AND current_x < (x"10E"+ DIGITLENGHT) AND current_y >=  FINALHIGH AND current_y < (FINALHIGH + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(milhar)(to_Integer(UNSIGNED(current_y- FINALHIGH)),to_Integer(UNSIGNED(current_x- x"10E"))));
            elsIF(current_x >= x"121" AND current_x < (x"121"+ DIGITLENGHT) AND current_y >=  FINALHIGH AND current_y < (FINALHIGH + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(centenas)(to_Integer(UNSIGNED(current_y- FINALHIGH)),to_Integer(UNSIGNED(current_x- x"121"))));
            elsIF(current_x >= x"134" AND current_x < (x"134"+ DIGITLENGHT) AND current_y >=  FINALHIGH AND current_y < (FINALHIGH + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(dezenas)(to_Integer(UNSIGNED(current_y- FINALHIGH)),to_Integer(UNSIGNED(current_x- x"134"))));
            elsIF(current_x >= x"147" AND current_x < (x"147"+ DIGITLENGHT) AND current_y >=  FINALHIGH AND current_y < (FINALHIGH + DIGITHIGH)) THEN
                colorOut(11 downto 8) <= (OTHERS => bcd_to_digit6x8(unidade)(to_Integer(UNSIGNED(current_y- FINALHIGH)),to_Integer(UNSIGNED(current_x- x"147"))));
            elsiF(counter(26)='0' and current_x >= x"D0" AND current_x < (x"D0"+ x"2E" ) AND current_y >=  x"7F" AND current_y < (x"7F" + x"E")) THEN
	            colorOut(11 downto 8) <= (OTHERS => Win(to_Integer(UNSIGNED(current_y- x"7F")),to_Integer(UNSIGNED(current_x- x"D0"))));   
	        elsiF(counter(26)='1' and current_x >= x"D0" AND current_x < (x"D0"+ x"2E" ) AND current_y >=  x"7F" AND current_y < (x"7F" + x"E")) THEN
	            colorOut(7 downto 4) <= (OTHERS => Win(to_Integer(UNSIGNED(current_y- x"7F")),to_Integer(UNSIGNED(current_x- x"D0"))));   
	        end if;    
        end if;
        
     end process;
        
end Behavioral;
